module top;

wire s;
initial
begin
    $display("hello");
    $finish;
end

endmodule
